// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

`timescale 1 ns / 1 ps

`include "uprj_netlists.v" // this file gets created automatically by multi_project_tools from the source section of info.yaml
`include "caravel_netlists.v"
`include "spiflash.v"

module zube_tb;
	initial begin
		$dumpfile ("zube.vcd");
		$dumpvars (0, zube_tb);
		#1;
	end

	reg clk;
	reg RSTB;
	reg power1, power2;
	reg power3, power4;

	wire gpio;
	wire [37:0] mprj_io;

	///// convenience signals that match what the cocotb test modules are looking for

	wire [7:0] z80_address_bus;
	wire [7:0] z80_data_bus_in;
	wire z80_write_strobe_b;
	wire z80_read_strobe_b;

	// 0-7 are management
	assign mprj_io[15:8] = z80_address_bus;
	// These are bidirectional
	assign mprj_io[23:16] = z80_data_bus_in;
	wire [7:0] z80_data_bus_out = mprj_io[23:16];
	assign mprj_io[24] = z80_write_strobe_b;
	assign mprj_io[25] = z80_read_strobe_b;
	wire z80_bus_dir = mprj_io[26];
	// 27 and higher are unused
	/////

	wire flash_csb;
	wire flash_clk;
	wire flash_io0;
	wire flash_io1;

	wire VDD3V3 = power1;
	wire VDD1V8 = power2;
	wire USER_VDD3V3 = power3;
	wire USER_VDD1V8 = power4;
	wire VSS = 1'b0;

	caravel uut(
		.vddio    (VDD3V3),
		.vssio    (VSS),
		.vdda     (VDD3V3),
		.vssa     (VSS),
		.vccd     (VDD1V8),
		.vssd     (VSS),
		.vdda1    (USER_VDD3V3),
		.vdda2    (USER_VDD3V3),
		.vssa1    (VSS),
		.vssa2    (VSS),
		.vccd1    (USER_VDD1V8),
		.vccd2    (USER_VDD1V8),
		.vssd1    (VSS),
		.vssd2    (VSS),
		.clock    (clk),
		.gpio     (gpio),
		.mprj_io  (mprj_io),
		.flash_csb(flash_csb),
		.flash_clk(flash_clk),
		.flash_io0(flash_io0),
		.flash_io1(flash_io1),
		.resetb   (RSTB)
	);

	spiflash #(
		.FILENAME("zube.hex")
	) spiflash (
		.csb(flash_csb),
		.clk(flash_clk),
		.io0(flash_io0),
		.io1(flash_io1),
		.io2(),          // not used
		.io3()           // not used
	);

endmodule
`default_nettype wire
